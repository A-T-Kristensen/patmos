library verilog;
use verilog.vl_types.all;
entity \InOut\ is
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        io_memInOut_M_Cmd: in     vl_logic_vector(2 downto 0);
        io_memInOut_M_Addr: in     vl_logic_vector(31 downto 0);
        io_memInOut_M_Data: in     vl_logic_vector(31 downto 0);
        io_memInOut_M_ByteEn: in     vl_logic_vector(3 downto 0);
        io_memInOut_S_Resp: out    vl_logic_vector(1 downto 0);
        io_memInOut_S_Data: out    vl_logic_vector(31 downto 0);
        io_comConf_M_Cmd: out    vl_logic_vector(2 downto 0);
        io_comConf_M_Addr: out    vl_logic_vector(31 downto 0);
        io_comConf_M_Data: out    vl_logic_vector(31 downto 0);
        io_comConf_M_ByteEn: out    vl_logic_vector(3 downto 0);
        io_comConf_M_RespAccept: out    vl_logic;
        io_comConf_S_Resp: in     vl_logic_vector(1 downto 0);
        io_comConf_S_Data: in     vl_logic_vector(31 downto 0);
        io_comConf_S_CmdAccept: in     vl_logic;
        io_comConf_S_Reset_n: in     vl_logic;
        io_comConf_S_Flag: in     vl_logic_vector(1 downto 0);
        io_comSpm_M_Cmd : out    vl_logic_vector(2 downto 0);
        io_comSpm_M_Addr: out    vl_logic_vector(31 downto 0);
        io_comSpm_M_Data: out    vl_logic_vector(31 downto 0);
        io_comSpm_M_ByteEn: out    vl_logic_vector(3 downto 0);
        io_comSpm_S_Resp: in     vl_logic_vector(1 downto 0);
        io_comSpm_S_Data: in     vl_logic_vector(31 downto 0);
        io_excInOut_M_Cmd: out    vl_logic_vector(2 downto 0);
        io_excInOut_M_Addr: out    vl_logic_vector(31 downto 0);
        io_excInOut_M_Data: out    vl_logic_vector(31 downto 0);
        io_excInOut_M_ByteEn: out    vl_logic_vector(3 downto 0);
        io_excInOut_S_Resp: in     vl_logic_vector(1 downto 0);
        io_excInOut_S_Data: in     vl_logic_vector(31 downto 0);
        io_intrs_15     : out    vl_logic;
        io_intrs_14     : out    vl_logic;
        io_intrs_13     : out    vl_logic;
        io_intrs_12     : out    vl_logic;
        io_intrs_11     : out    vl_logic;
        io_intrs_10     : out    vl_logic;
        io_intrs_9      : out    vl_logic;
        io_intrs_8      : out    vl_logic;
        io_intrs_7      : out    vl_logic;
        io_intrs_6      : out    vl_logic;
        io_intrs_5      : out    vl_logic;
        io_intrs_4      : out    vl_logic;
        io_intrs_3      : out    vl_logic;
        io_intrs_2      : out    vl_logic;
        io_intrs_1      : out    vl_logic;
        io_intrs_0      : out    vl_logic;
        io_superMode    : in     vl_logic;
        io_internalIO_perf_ic_hit: in     vl_logic;
        io_internalIO_perf_ic_miss: in     vl_logic;
        io_internalIO_perf_dc_hit: in     vl_logic;
        io_internalIO_perf_dc_miss: in     vl_logic;
        io_internalIO_perf_sc_spill: in     vl_logic;
        io_internalIO_perf_sc_fill: in     vl_logic;
        io_internalIO_perf_wc_hit: in     vl_logic;
        io_internalIO_perf_wc_miss: in     vl_logic;
        io_internalIO_perf_mem_read: in     vl_logic;
        io_internalIO_perf_mem_write: in     vl_logic;
        io_uartPins_tx  : out    vl_logic;
        io_uartPins_rx  : in     vl_logic;
        io_ledsPins_led : out    vl_logic_vector(8 downto 0);
        io_keysPins_key : in     vl_logic_vector(3 downto 0);
        io_cpuInfoPins_id: in     vl_logic_vector(31 downto 0);
        io_cpuInfoPins_cnt: in     vl_logic_vector(31 downto 0)
    );
end \InOut\;
